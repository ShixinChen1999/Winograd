module Transfer( // @[:@81.2]
  input        clock, // @[:@82.4]
  input        reset, // @[:@83.4]
  input  [7:0] io_dIn, // @[:@84.4]
  input  [9:0] io_dIn_addr, // @[:@84.4]
  input        io_input_valid, // @[:@84.4]
  output [7:0] io_RAM_OUT_0, // @[:@84.4]
  output [7:0] io_RAM_OUT_1, // @[:@84.4]
  output [7:0] io_RAM_OUT_2, // @[:@84.4]
  output [7:0] io_RAM_OUT_3, // @[:@84.4]
  output [7:0] io_RAM_OUT_4, // @[:@84.4]
  output [7:0] io_RAM_OUT_5, // @[:@84.4]
  output       io_out_valid // @[:@84.4]
);
  wire [15:0] DualPortRAM_io_dataOut; // @[transfer.scala 93:39:@97.4]
  wire  DualPortRAM_io_output_valid; // @[transfer.scala 93:39:@97.4]
  wire [9:0] DualPortRAM_io_output_addr; // @[transfer.scala 93:39:@97.4]
  wire  DualPortRAM_io_input_valid; // @[transfer.scala 93:39:@97.4]
  wire [15:0] DualPortRAM_io_dataIn; // @[transfer.scala 93:39:@97.4]
  wire [9:0] DualPortRAM_io_in_addr; // @[transfer.scala 93:39:@97.4]
  wire  DualPortRAM_reset; // @[transfer.scala 93:39:@97.4]
  wire  DualPortRAM_clock; // @[transfer.scala 93:39:@97.4]
  wire [15:0] DualPortRAM_1_io_dataOut; // @[transfer.scala 93:39:@106.4]
  wire  DualPortRAM_1_io_output_valid; // @[transfer.scala 93:39:@106.4]
  wire [9:0] DualPortRAM_1_io_output_addr; // @[transfer.scala 93:39:@106.4]
  wire  DualPortRAM_1_io_input_valid; // @[transfer.scala 93:39:@106.4]
  wire [15:0] DualPortRAM_1_io_dataIn; // @[transfer.scala 93:39:@106.4]
  wire [9:0] DualPortRAM_1_io_in_addr; // @[transfer.scala 93:39:@106.4]
  wire  DualPortRAM_1_reset; // @[transfer.scala 93:39:@106.4]
  wire  DualPortRAM_1_clock; // @[transfer.scala 93:39:@106.4]
  wire [15:0] DualPortRAM_2_io_dataOut; // @[transfer.scala 93:39:@115.4]
  wire  DualPortRAM_2_io_output_valid; // @[transfer.scala 93:39:@115.4]
  wire [9:0] DualPortRAM_2_io_output_addr; // @[transfer.scala 93:39:@115.4]
  wire  DualPortRAM_2_io_input_valid; // @[transfer.scala 93:39:@115.4]
  wire [15:0] DualPortRAM_2_io_dataIn; // @[transfer.scala 93:39:@115.4]
  wire [9:0] DualPortRAM_2_io_in_addr; // @[transfer.scala 93:39:@115.4]
  wire  DualPortRAM_2_reset; // @[transfer.scala 93:39:@115.4]
  wire  DualPortRAM_2_clock; // @[transfer.scala 93:39:@115.4]
  wire [15:0] DualPortRAM_3_io_dataOut; // @[transfer.scala 93:39:@124.4]
  wire  DualPortRAM_3_io_output_valid; // @[transfer.scala 93:39:@124.4]
  wire [9:0] DualPortRAM_3_io_output_addr; // @[transfer.scala 93:39:@124.4]
  wire  DualPortRAM_3_io_input_valid; // @[transfer.scala 93:39:@124.4]
  wire [15:0] DualPortRAM_3_io_dataIn; // @[transfer.scala 93:39:@124.4]
  wire [9:0] DualPortRAM_3_io_in_addr; // @[transfer.scala 93:39:@124.4]
  wire  DualPortRAM_3_reset; // @[transfer.scala 93:39:@124.4]
  wire  DualPortRAM_3_clock; // @[transfer.scala 93:39:@124.4]
  wire [15:0] DualPortRAM_4_io_dataOut; // @[transfer.scala 93:39:@133.4]
  wire  DualPortRAM_4_io_output_valid; // @[transfer.scala 93:39:@133.4]
  wire [9:0] DualPortRAM_4_io_output_addr; // @[transfer.scala 93:39:@133.4]
  wire  DualPortRAM_4_io_input_valid; // @[transfer.scala 93:39:@133.4]
  wire [15:0] DualPortRAM_4_io_dataIn; // @[transfer.scala 93:39:@133.4]
  wire [9:0] DualPortRAM_4_io_in_addr; // @[transfer.scala 93:39:@133.4]
  wire  DualPortRAM_4_reset; // @[transfer.scala 93:39:@133.4]
  wire  DualPortRAM_4_clock; // @[transfer.scala 93:39:@133.4]
  wire [15:0] DualPortRAM_5_io_dataOut; // @[transfer.scala 93:39:@142.4]
  wire  DualPortRAM_5_io_output_valid; // @[transfer.scala 93:39:@142.4]
  wire [9:0] DualPortRAM_5_io_output_addr; // @[transfer.scala 93:39:@142.4]
  wire  DualPortRAM_5_io_input_valid; // @[transfer.scala 93:39:@142.4]
  wire [15:0] DualPortRAM_5_io_dataIn; // @[transfer.scala 93:39:@142.4]
  wire [9:0] DualPortRAM_5_io_in_addr; // @[transfer.scala 93:39:@142.4]
  wire  DualPortRAM_5_reset; // @[transfer.scala 93:39:@142.4]
  wire  DualPortRAM_5_clock; // @[transfer.scala 93:39:@142.4]
  reg [7:0] value; // @[Counter.scala 26:33:@86.4]
  reg [31:0] _RAND_0;
  wire  _T_38; // @[Counter.scala 34:24:@88.6]
  wire [8:0] _T_40; // @[Counter.scala 35:22:@89.6]
  wire [7:0] _T_41; // @[Counter.scala 35:22:@90.6]
  wire [7:0] _GEN_0; // @[Counter.scala 37:21:@92.6]
  wire [7:0] _GEN_1; // @[Counter.scala 63:17:@87.4]
  wire [7:0] _T_231; // @[transfer.scala 96:19:@200.4]
  wire [7:0] _GEN_2; // @[transfer.scala 96:31:@201.4]
  wire [2:0] NUM_RAM; // @[transfer.scala 96:31:@201.4]
  wire  _T_238; // @[transfer.scala 99:28:@204.4]
  wire  _T_244; // @[transfer.scala 99:56:@207.4]
  wire  _T_245; // @[transfer.scala 99:34:@208.4]
  wire [7:0] _GEN_3; // @[transfer.scala 100:26:@211.6]
  wire [1:0] _T_249; // @[transfer.scala 100:26:@211.6]
  wire  _T_251; // @[transfer.scala 100:30:@212.6]
  wire [7:0] _GEN_4; // @[transfer.scala 100:41:@213.6]
  wire [1:0] _T_253; // @[transfer.scala 100:41:@213.6]
  wire  _T_255; // @[transfer.scala 100:45:@214.6]
  wire  _T_256; // @[transfer.scala 100:36:@215.6]
  wire [9:0] _GEN_5; // @[transfer.scala 101:37:@217.8]
  wire [4:0] _T_258; // @[transfer.scala 101:37:@217.8]
  wire  _T_279; // @[transfer.scala 107:51:@272.8]
  wire  _T_280; // @[transfer.scala 107:42:@273.8]
  wire  _T_299; // @[transfer.scala 114:36:@328.10]
  wire  _T_304; // @[transfer.scala 114:42:@331.10]
  wire  _GEN_8; // @[transfer.scala 114:58:@332.10]
  wire  _GEN_15; // @[transfer.scala 107:58:@274.8]
  wire [4:0] _GEN_16; // @[transfer.scala 107:58:@274.8]
  wire  _GEN_19; // @[transfer.scala 107:58:@274.8]
  wire  _GEN_26; // @[transfer.scala 100:52:@216.6]
  wire [4:0] _GEN_27; // @[transfer.scala 100:52:@216.6]
  wire  _GEN_30; // @[transfer.scala 100:52:@216.6]
  wire  _T_336; // @[transfer.scala 129:34:@438.6]
  wire  _T_342; // @[transfer.scala 129:62:@441.6]
  wire  _T_343; // @[transfer.scala 129:40:@442.6]
  wire  _GEN_103; // @[transfer.scala 129:69:@443.6]
  wire  _GEN_107; // @[transfer.scala 129:69:@443.6]
  wire  _GEN_112; // @[transfer.scala 129:69:@443.6]
  wire  _GEN_116; // @[transfer.scala 129:69:@443.6]
  reg  _T_516; // @[Reg.scala 11:16:@895.4]
  reg [31:0] _RAND_1;
  reg  _T_518; // @[Reg.scala 11:16:@899.4]
  reg [31:0] _RAND_2;
  reg  _T_520; // @[Reg.scala 11:16:@903.4]
  reg [31:0] _RAND_3;
  reg  _T_522; // @[Reg.scala 11:16:@907.4]
  reg [31:0] _RAND_4;
  reg  _T_524; // @[Reg.scala 11:16:@911.4]
  reg [31:0] _RAND_5;
  reg  _T_526; // @[Reg.scala 11:16:@915.4]
  reg [31:0] _RAND_6;
  reg  _T_528; // @[Reg.scala 11:16:@919.4]
  reg [31:0] _RAND_7;
  reg  _T_530; // @[Reg.scala 11:16:@923.4]
  reg [31:0] _RAND_8;
  reg  _T_532; // @[Reg.scala 11:16:@927.4]
  reg [31:0] _RAND_9;
  reg  _T_534; // @[Reg.scala 11:16:@931.4]
  reg [31:0] _RAND_10;
  reg  _T_536; // @[Reg.scala 11:16:@935.4]
  reg [31:0] _RAND_11;
  reg  _T_538; // @[Reg.scala 11:16:@939.4]
  reg [31:0] _RAND_12;
  reg  _T_540; // @[Reg.scala 11:16:@943.4]
  reg [31:0] _RAND_13;
  reg  _T_542; // @[Reg.scala 11:16:@947.4]
  reg [31:0] _RAND_14;
  reg  _T_544; // @[Reg.scala 11:16:@951.4]
  reg [31:0] _RAND_15;
  reg  _T_546; // @[Reg.scala 11:16:@955.4]
  reg [31:0] _RAND_16;
  reg  _T_548; // @[Reg.scala 11:16:@959.4]
  reg [31:0] _RAND_17;
  reg  _T_550; // @[Reg.scala 11:16:@963.4]
  reg [31:0] _RAND_18;
  reg  _T_552; // @[Reg.scala 11:16:@967.4]
  reg [31:0] _RAND_19;
  reg  _T_554; // @[Reg.scala 11:16:@971.4]
  reg [31:0] _RAND_20;
  reg  _T_556; // @[Reg.scala 11:16:@975.4]
  reg [31:0] _RAND_21;
  reg  _T_558; // @[Reg.scala 11:16:@979.4]
  reg [31:0] _RAND_22;
  reg  _T_560; // @[Reg.scala 11:16:@983.4]
  reg [31:0] _RAND_23;
  reg  _T_562; // @[Reg.scala 11:16:@987.4]
  reg [31:0] _RAND_24;
  reg  _T_564; // @[Reg.scala 11:16:@991.4]
  reg [31:0] _RAND_25;
  reg  _T_566; // @[Reg.scala 11:16:@995.4]
  reg [31:0] _RAND_26;
  reg  _T_568; // @[Reg.scala 11:16:@999.4]
  reg [31:0] _RAND_27;
  reg  _T_570; // @[Reg.scala 11:16:@1003.4]
  reg [31:0] _RAND_28;
  reg  _T_572; // @[Reg.scala 11:16:@1007.4]
  reg [31:0] _RAND_29;
  reg  _T_574; // @[Reg.scala 11:16:@1011.4]
  reg [31:0] _RAND_30;
  reg  _T_576; // @[Reg.scala 11:16:@1015.4]
  reg [31:0] _RAND_31;
  reg  _T_578; // @[Reg.scala 11:16:@1019.4]
  reg [31:0] _RAND_32;
  reg  _T_580; // @[Reg.scala 11:16:@1023.4]
  reg [31:0] _RAND_33;
  reg  _T_582; // @[Reg.scala 11:16:@1027.4]
  reg [31:0] _RAND_34;
  reg  _T_584; // @[Reg.scala 11:16:@1031.4]
  reg [31:0] _RAND_35;
  reg  _T_586; // @[Reg.scala 11:16:@1035.4]
  reg [31:0] _RAND_36;
  reg  _T_588; // @[Reg.scala 11:16:@1039.4]
  reg [31:0] _RAND_37;
  reg  _T_590; // @[Reg.scala 11:16:@1043.4]
  reg [31:0] _RAND_38;
  reg  _T_592; // @[Reg.scala 11:16:@1047.4]
  reg [31:0] _RAND_39;
  reg  _T_594; // @[Reg.scala 11:16:@1051.4]
  reg [31:0] _RAND_40;
  reg  _T_596; // @[Reg.scala 11:16:@1055.4]
  reg [31:0] _RAND_41;
  reg  _T_598; // @[Reg.scala 11:16:@1059.4]
  reg [31:0] _RAND_42;
  reg  _T_600; // @[Reg.scala 11:16:@1063.4]
  reg [31:0] _RAND_43;
  reg  _T_602; // @[Reg.scala 11:16:@1067.4]
  reg [31:0] _RAND_44;
  reg  _T_604; // @[Reg.scala 11:16:@1071.4]
  reg [31:0] _RAND_45;
  reg  _T_606; // @[Reg.scala 11:16:@1075.4]
  reg [31:0] _RAND_46;
  reg  _T_608; // @[Reg.scala 11:16:@1079.4]
  reg [31:0] _RAND_47;
  reg  _T_610; // @[Reg.scala 11:16:@1083.4]
  reg [31:0] _RAND_48;
  reg  _T_612; // @[Reg.scala 11:16:@1087.4]
  reg [31:0] _RAND_49;
  reg  _T_614; // @[Reg.scala 11:16:@1091.4]
  reg [31:0] _RAND_50;
  reg  _T_616; // @[Reg.scala 11:16:@1095.4]
  reg [31:0] _RAND_51;
  reg  _T_618; // @[Reg.scala 11:16:@1099.4]
  reg [31:0] _RAND_52;
  reg  _T_620; // @[Reg.scala 11:16:@1103.4]
  reg [31:0] _RAND_53;
  reg  _T_622; // @[Reg.scala 11:16:@1107.4]
  reg [31:0] _RAND_54;
  reg  _T_624; // @[Reg.scala 11:16:@1111.4]
  reg [31:0] _RAND_55;
  reg  _T_626; // @[Reg.scala 11:16:@1115.4]
  reg [31:0] _RAND_56;
  reg  _T_628; // @[Reg.scala 11:16:@1119.4]
  reg [31:0] _RAND_57;
  reg  _T_630; // @[Reg.scala 11:16:@1123.4]
  reg [31:0] _RAND_58;
  reg  _T_632; // @[Reg.scala 11:16:@1127.4]
  reg [31:0] _RAND_59;
  reg  _T_634; // @[Reg.scala 11:16:@1131.4]
  reg [31:0] _RAND_60;
  reg  _T_636; // @[Reg.scala 11:16:@1135.4]
  reg [31:0] _RAND_61;
  reg  _T_638; // @[Reg.scala 11:16:@1139.4]
  reg [31:0] _RAND_62;
  reg  _T_640; // @[Reg.scala 11:16:@1143.4]
  reg [31:0] _RAND_63;
  reg  _T_642; // @[Reg.scala 11:16:@1147.4]
  reg [31:0] _RAND_64;
  reg [7:0] value_1; // @[Counter.scala 26:33:@1152.4]
  reg [31:0] _RAND_65;
  wire  _T_646; // @[Counter.scala 34:24:@1154.6]
  wire [8:0] _T_648; // @[Counter.scala 35:22:@1155.6]
  wire [7:0] _T_649; // @[Counter.scala 35:22:@1156.6]
  wire [7:0] _GEN_210; // @[Counter.scala 37:21:@1158.6]
  wire [7:0] _GEN_211; // @[Counter.scala 63:17:@1153.4]
  wire [7:0] dOut_addr; // @[transfer.scala 195:24:@1163.4]
  wire [7:0] _GEN_6; // @[transfer.scala 199:17:@1170.6]
  wire [1:0] _T_666; // @[transfer.scala 199:17:@1170.6]
  wire  _T_668; // @[transfer.scala 199:21:@1171.6]
  wire [7:0] _T_670; // @[transfer.scala 200:20:@1173.8]
  wire [7:0] _GEN_7; // @[transfer.scala 200:32:@1174.8]
  wire [2:0] _T_672; // @[transfer.scala 200:32:@1174.8]
  wire  _T_674; // @[transfer.scala 200:36:@1175.8]
  wire  _T_680; // @[transfer.scala 200:68:@1178.8]
  wire  _T_681; // @[transfer.scala 200:42:@1179.8]
  wire [7:0] _GEN_9; // @[transfer.scala 201:34:@1182.10]
  wire [2:0] _T_685; // @[transfer.scala 201:34:@1182.10]
  wire  _T_687; // @[transfer.scala 201:38:@1183.10]
  wire [7:0] _GEN_10; // @[transfer.scala 202:51:@1185.12]
  wire [4:0] _T_689; // @[transfer.scala 202:51:@1185.12]
  wire [4:0] _GEN_215; // @[transfer.scala 201:45:@1184.10]
  wire  _T_717; // @[transfer.scala 212:42:@1264.10]
  wire  _T_723; // @[transfer.scala 212:74:@1267.10]
  wire  _T_724; // @[transfer.scala 212:48:@1268.10]
  wire  _T_760; // @[transfer.scala 224:42:@1353.12]
  wire  _T_766; // @[transfer.scala 224:74:@1356.12]
  wire  _T_767; // @[transfer.scala 224:48:@1357.12]
  wire  _GEN_290; // @[transfer.scala 212:81:@1269.10]
  wire [4:0] _GEN_291; // @[transfer.scala 212:81:@1269.10]
  wire  _GEN_304; // @[transfer.scala 212:81:@1269.10]
  wire  _GEN_316; // @[transfer.scala 200:75:@1180.8]
  wire [4:0] _GEN_317; // @[transfer.scala 200:75:@1180.8]
  wire  _GEN_330; // @[transfer.scala 200:75:@1180.8]
  wire  _GEN_344; // @[transfer.scala 200:75:@1180.8]
  wire  _GEN_356; // @[transfer.scala 199:28:@1172.6]
  wire  _GEN_370; // @[transfer.scala 199:28:@1172.6]
  wire  _GEN_384; // @[transfer.scala 199:28:@1172.6]
  DualPortRAM DualPortRAM ( // @[transfer.scala 93:39:@97.4]
    .io_dataOut(DualPortRAM_io_dataOut),
    .io_output_valid(DualPortRAM_io_output_valid),
    .io_output_addr(DualPortRAM_io_output_addr),
    .io_input_valid(DualPortRAM_io_input_valid),
    .io_dataIn(DualPortRAM_io_dataIn),
    .io_in_addr(DualPortRAM_io_in_addr),
    .reset(DualPortRAM_reset),
    .clock(DualPortRAM_clock)
  );
  DualPortRAM DualPortRAM_1 ( // @[transfer.scala 93:39:@106.4]
    .io_dataOut(DualPortRAM_1_io_dataOut),
    .io_output_valid(DualPortRAM_1_io_output_valid),
    .io_output_addr(DualPortRAM_1_io_output_addr),
    .io_input_valid(DualPortRAM_1_io_input_valid),
    .io_dataIn(DualPortRAM_1_io_dataIn),
    .io_in_addr(DualPortRAM_1_io_in_addr),
    .reset(DualPortRAM_1_reset),
    .clock(DualPortRAM_1_clock)
  );
  DualPortRAM DualPortRAM_2 ( // @[transfer.scala 93:39:@115.4]
    .io_dataOut(DualPortRAM_2_io_dataOut),
    .io_output_valid(DualPortRAM_2_io_output_valid),
    .io_output_addr(DualPortRAM_2_io_output_addr),
    .io_input_valid(DualPortRAM_2_io_input_valid),
    .io_dataIn(DualPortRAM_2_io_dataIn),
    .io_in_addr(DualPortRAM_2_io_in_addr),
    .reset(DualPortRAM_2_reset),
    .clock(DualPortRAM_2_clock)
  );
  DualPortRAM DualPortRAM_3 ( // @[transfer.scala 93:39:@124.4]
    .io_dataOut(DualPortRAM_3_io_dataOut),
    .io_output_valid(DualPortRAM_3_io_output_valid),
    .io_output_addr(DualPortRAM_3_io_output_addr),
    .io_input_valid(DualPortRAM_3_io_input_valid),
    .io_dataIn(DualPortRAM_3_io_dataIn),
    .io_in_addr(DualPortRAM_3_io_in_addr),
    .reset(DualPortRAM_3_reset),
    .clock(DualPortRAM_3_clock)
  );
  DualPortRAM DualPortRAM_4 ( // @[transfer.scala 93:39:@133.4]
    .io_dataOut(DualPortRAM_4_io_dataOut),
    .io_output_valid(DualPortRAM_4_io_output_valid),
    .io_output_addr(DualPortRAM_4_io_output_addr),
    .io_input_valid(DualPortRAM_4_io_input_valid),
    .io_dataIn(DualPortRAM_4_io_dataIn),
    .io_in_addr(DualPortRAM_4_io_in_addr),
    .reset(DualPortRAM_4_reset),
    .clock(DualPortRAM_4_clock)
  );
  DualPortRAM DualPortRAM_5 ( // @[transfer.scala 93:39:@142.4]
    .io_dataOut(DualPortRAM_5_io_dataOut),
    .io_output_valid(DualPortRAM_5_io_output_valid),
    .io_output_addr(DualPortRAM_5_io_output_addr),
    .io_input_valid(DualPortRAM_5_io_input_valid),
    .io_dataIn(DualPortRAM_5_io_dataIn),
    .io_in_addr(DualPortRAM_5_io_in_addr),
    .reset(DualPortRAM_5_reset),
    .clock(DualPortRAM_5_clock)
  );
  assign _T_38 = value == 8'hbf; // @[Counter.scala 34:24:@88.6]
  assign _T_40 = value + 8'h1; // @[Counter.scala 35:22:@89.6]
  assign _T_41 = _T_40[7:0]; // @[Counter.scala 35:22:@90.6]
  assign _GEN_0 = _T_38 ? 8'h0 : _T_41; // @[Counter.scala 37:21:@92.6]
  assign _GEN_1 = io_input_valid ? _GEN_0 : value; // @[Counter.scala 63:17:@87.4]
  assign _T_231 = value / 8'h10; // @[transfer.scala 96:19:@200.4]
  assign _GEN_2 = _T_231 % 8'h6; // @[transfer.scala 96:31:@201.4]
  assign NUM_RAM = _GEN_2[2:0]; // @[transfer.scala 96:31:@201.4]
  assign _T_238 = NUM_RAM == 3'h0; // @[transfer.scala 99:28:@204.4]
  assign _T_244 = NUM_RAM == 3'h1; // @[transfer.scala 99:56:@207.4]
  assign _T_245 = _T_238 | _T_244; // @[transfer.scala 99:34:@208.4]
  assign _GEN_3 = _T_231 % 8'h2; // @[transfer.scala 100:26:@211.6]
  assign _T_249 = _GEN_3[1:0]; // @[transfer.scala 100:26:@211.6]
  assign _T_251 = _T_249 == 2'h0; // @[transfer.scala 100:30:@212.6]
  assign _GEN_4 = value % 8'h2; // @[transfer.scala 100:41:@213.6]
  assign _T_253 = _GEN_4[1:0]; // @[transfer.scala 100:41:@213.6]
  assign _T_255 = _T_253 == 2'h0; // @[transfer.scala 100:45:@214.6]
  assign _T_256 = _T_251 & _T_255; // @[transfer.scala 100:36:@215.6]
  assign _GEN_5 = io_dIn_addr % 10'h10; // @[transfer.scala 101:37:@217.8]
  assign _T_258 = _GEN_5[4:0]; // @[transfer.scala 101:37:@217.8]
  assign _T_279 = _T_253 == 2'h1; // @[transfer.scala 107:51:@272.8]
  assign _T_280 = _T_251 & _T_279; // @[transfer.scala 107:42:@273.8]
  assign _T_299 = _T_249 == 2'h1; // @[transfer.scala 114:36:@328.10]
  assign _T_304 = _T_299 & _T_255; // @[transfer.scala 114:42:@331.10]
  assign _GEN_8 = _T_304 ? 1'h0 : 1'h1; // @[transfer.scala 114:58:@332.10]
  assign _GEN_15 = _T_280 ? 1'h1 : _T_304; // @[transfer.scala 107:58:@274.8]
  assign _GEN_16 = _T_280 ? _T_258 : _T_258; // @[transfer.scala 107:58:@274.8]
  assign _GEN_19 = _T_280 ? 1'h0 : _GEN_8; // @[transfer.scala 107:58:@274.8]
  assign _GEN_26 = _T_256 ? 1'h1 : _GEN_19; // @[transfer.scala 100:52:@216.6]
  assign _GEN_27 = _T_256 ? _T_258 : _T_258; // @[transfer.scala 100:52:@216.6]
  assign _GEN_30 = _T_256 ? 1'h0 : _GEN_15; // @[transfer.scala 100:52:@216.6]
  assign _T_336 = NUM_RAM == 3'h2; // @[transfer.scala 129:34:@438.6]
  assign _T_342 = NUM_RAM == 3'h3; // @[transfer.scala 129:62:@441.6]
  assign _T_343 = _T_336 | _T_342; // @[transfer.scala 129:40:@442.6]
  assign _GEN_103 = _T_343 ? _GEN_26 : 1'h0; // @[transfer.scala 129:69:@443.6]
  assign _GEN_107 = _T_343 ? _GEN_30 : 1'h0; // @[transfer.scala 129:69:@443.6]
  assign _GEN_112 = _T_343 ? 1'h0 : _GEN_26; // @[transfer.scala 129:69:@443.6]
  assign _GEN_116 = _T_343 ? 1'h0 : _GEN_30; // @[transfer.scala 129:69:@443.6]
  assign _T_646 = value_1 == 8'hbf; // @[Counter.scala 34:24:@1154.6]
  assign _T_648 = value_1 + 8'h1; // @[Counter.scala 35:22:@1155.6]
  assign _T_649 = _T_648[7:0]; // @[Counter.scala 35:22:@1156.6]
  assign _GEN_210 = _T_646 ? 8'h0 : _T_649; // @[Counter.scala 37:21:@1158.6]
  assign _GEN_211 = io_out_valid ? _GEN_210 : value_1; // @[Counter.scala 63:17:@1153.4]
  assign dOut_addr = value_1 / 8'h2; // @[transfer.scala 195:24:@1163.4]
  assign _GEN_6 = value_1 % 8'h2; // @[transfer.scala 199:17:@1170.6]
  assign _T_666 = _GEN_6[1:0]; // @[transfer.scala 199:17:@1170.6]
  assign _T_668 = _T_666 == 2'h0; // @[transfer.scala 199:21:@1171.6]
  assign _T_670 = value_1 / 8'h10; // @[transfer.scala 200:20:@1173.8]
  assign _GEN_7 = _T_670 % 8'h6; // @[transfer.scala 200:32:@1174.8]
  assign _T_672 = _GEN_7[2:0]; // @[transfer.scala 200:32:@1174.8]
  assign _T_674 = _T_672 == 3'h0; // @[transfer.scala 200:36:@1175.8]
  assign _T_680 = _T_672 == 3'h1; // @[transfer.scala 200:68:@1178.8]
  assign _T_681 = _T_674 | _T_680; // @[transfer.scala 200:42:@1179.8]
  assign _GEN_9 = _T_670 % 8'h4; // @[transfer.scala 201:34:@1182.10]
  assign _T_685 = _GEN_9[2:0]; // @[transfer.scala 201:34:@1182.10]
  assign _T_687 = _T_685 == 3'h0; // @[transfer.scala 201:38:@1183.10]
  assign _GEN_10 = dOut_addr % 8'h10; // @[transfer.scala 202:51:@1185.12]
  assign _T_689 = _GEN_10[4:0]; // @[transfer.scala 202:51:@1185.12]
  assign _GEN_215 = _T_687 ? _T_689 : _T_689; // @[transfer.scala 201:45:@1184.10]
  assign _T_717 = _T_672 == 3'h2; // @[transfer.scala 212:42:@1264.10]
  assign _T_723 = _T_672 == 3'h3; // @[transfer.scala 212:74:@1267.10]
  assign _T_724 = _T_717 | _T_723; // @[transfer.scala 212:48:@1268.10]
  assign _T_760 = _T_672 == 3'h4; // @[transfer.scala 224:42:@1353.12]
  assign _T_766 = _T_672 == 3'h5; // @[transfer.scala 224:74:@1356.12]
  assign _T_767 = _T_760 | _T_766; // @[transfer.scala 224:48:@1357.12]
  assign _GEN_290 = _T_724 ? 1'h1 : _T_767; // @[transfer.scala 212:81:@1269.10]
  assign _GEN_291 = _T_724 ? _GEN_215 : _GEN_215; // @[transfer.scala 212:81:@1269.10]
  assign _GEN_304 = _T_724 ? 1'h0 : _T_767; // @[transfer.scala 212:81:@1269.10]
  assign _GEN_316 = _T_681 ? 1'h1 : _GEN_304; // @[transfer.scala 200:75:@1180.8]
  assign _GEN_317 = _T_681 ? _GEN_215 : _GEN_215; // @[transfer.scala 200:75:@1180.8]
  assign _GEN_330 = _T_681 ? 1'h1 : _T_724; // @[transfer.scala 200:75:@1180.8]
  assign _GEN_344 = _T_681 ? 1'h0 : _GEN_290; // @[transfer.scala 200:75:@1180.8]
  assign _GEN_356 = _T_668 ? _GEN_316 : 1'h0; // @[transfer.scala 199:28:@1172.6]
  assign _GEN_370 = _T_668 ? _GEN_330 : 1'h0; // @[transfer.scala 199:28:@1172.6]
  assign _GEN_384 = _T_668 ? _GEN_344 : 1'h0; // @[transfer.scala 199:28:@1172.6]
   assign io_RAM_OUT_0 = DualPortRAM_io_dataOut;
           assign io_RAM_OUT_1 = DualPortRAM_1_io_dataOut;
           assign io_RAM_OUT_2 =  DualPortRAM_2_io_dataOut;
           assign io_RAM_OUT_3 =  DualPortRAM_3_io_dataOut;
           assign io_RAM_OUT_4 =  DualPortRAM_4_io_dataOut;
           assign io_RAM_OUT_5 =  DualPortRAM_5_io_dataOut;
  assign io_out_valid = _T_642; // @[transfer.scala 191:15:@1151.4]
  assign DualPortRAM_io_output_valid = io_out_valid ? _GEN_356 : 1'h0; // @[transfer.scala 93:20:@153.4]
  assign DualPortRAM_io_output_addr = {{5'd0}, _GEN_317}; // @[transfer.scala 93:20:@154.4]
  assign DualPortRAM_io_input_valid = _T_245 ? _GEN_26 : 1'h0; // @[transfer.scala 93:20:@155.4]
  assign DualPortRAM_io_dataIn = {{8'd0}, io_dIn}; // @[transfer.scala 93:20:@156.4]
  assign DualPortRAM_io_in_addr = {{5'd0}, _GEN_27}; // @[transfer.scala 93:20:@157.4]
  assign DualPortRAM_reset = reset; // @[transfer.scala 93:20:@158.4]
  assign DualPortRAM_clock = clock; // @[transfer.scala 93:20:@159.4]
  assign DualPortRAM_1_io_output_valid = io_out_valid ? _GEN_356 : 1'h0; // @[transfer.scala 93:20:@161.4]
  assign DualPortRAM_1_io_output_addr = {{5'd0}, _GEN_317}; // @[transfer.scala 93:20:@162.4]
  assign DualPortRAM_1_io_input_valid = _T_245 ? _GEN_30 : 1'h0; // @[transfer.scala 93:20:@163.4]
  assign DualPortRAM_1_io_dataIn = {{8'd0}, io_dIn}; // @[transfer.scala 93:20:@164.4]
  assign DualPortRAM_1_io_in_addr = {{5'd0}, _GEN_16}; // @[transfer.scala 93:20:@165.4]
  assign DualPortRAM_1_reset = reset; // @[transfer.scala 93:20:@166.4]
  assign DualPortRAM_1_clock = clock; // @[transfer.scala 93:20:@167.4]
  assign DualPortRAM_2_io_output_valid = io_out_valid ? _GEN_370 : 1'h0; // @[transfer.scala 93:20:@169.4]
  assign DualPortRAM_2_io_output_addr = {{5'd0}, _GEN_317}; // @[transfer.scala 93:20:@170.4]
  assign DualPortRAM_2_io_input_valid = _T_245 ? 1'h0 : _GEN_103; // @[transfer.scala 93:20:@171.4]
  assign DualPortRAM_2_io_dataIn = {{8'd0}, io_dIn}; // @[transfer.scala 93:20:@172.4]
  assign DualPortRAM_2_io_in_addr = {{5'd0}, _GEN_27}; // @[transfer.scala 93:20:@173.4]
  assign DualPortRAM_2_reset = reset; // @[transfer.scala 93:20:@174.4]
  assign DualPortRAM_2_clock = clock; // @[transfer.scala 93:20:@175.4]
  assign DualPortRAM_3_io_output_valid = io_out_valid ? _GEN_370 : 1'h0; // @[transfer.scala 93:20:@177.4]
  assign DualPortRAM_3_io_output_addr = {{5'd0}, _GEN_317}; // @[transfer.scala 93:20:@178.4]
  assign DualPortRAM_3_io_input_valid = _T_245 ? 1'h0 : _GEN_107; // @[transfer.scala 93:20:@179.4]
  assign DualPortRAM_3_io_dataIn = {{8'd0}, io_dIn}; // @[transfer.scala 93:20:@180.4]
  assign DualPortRAM_3_io_in_addr = {{5'd0}, _GEN_16}; // @[transfer.scala 93:20:@181.4]
  assign DualPortRAM_3_reset = reset; // @[transfer.scala 93:20:@182.4]
  assign DualPortRAM_3_clock = clock; // @[transfer.scala 93:20:@183.4]
  assign DualPortRAM_4_io_output_valid = io_out_valid ? _GEN_384 : 1'h0; // @[transfer.scala 93:20:@185.4]
  assign DualPortRAM_4_io_output_addr = {{5'd0}, _GEN_291}; // @[transfer.scala 93:20:@186.4]
  assign DualPortRAM_4_io_input_valid = _T_245 ? 1'h0 : _GEN_112; // @[transfer.scala 93:20:@187.4]
  assign DualPortRAM_4_io_dataIn = {{8'd0}, io_dIn}; // @[transfer.scala 93:20:@188.4]
  assign DualPortRAM_4_io_in_addr = {{5'd0}, _GEN_27}; // @[transfer.scala 93:20:@189.4]
  assign DualPortRAM_4_reset = reset; // @[transfer.scala 93:20:@190.4]
  assign DualPortRAM_4_clock = clock; // @[transfer.scala 93:20:@191.4]
  assign DualPortRAM_5_io_output_valid = io_out_valid ? _GEN_384 : 1'h0; // @[transfer.scala 93:20:@193.4]
  assign DualPortRAM_5_io_output_addr = {{5'd0}, _GEN_291}; // @[transfer.scala 93:20:@194.4]
  assign DualPortRAM_5_io_input_valid = _T_245 ? 1'h0 : _GEN_116; // @[transfer.scala 93:20:@195.4]
  assign DualPortRAM_5_io_dataIn = {{8'd0}, io_dIn}; // @[transfer.scala 93:20:@196.4]
  assign DualPortRAM_5_io_in_addr = {{5'd0}, _GEN_16}; // @[transfer.scala 93:20:@197.4]
  assign DualPortRAM_5_reset = reset; // @[transfer.scala 93:20:@198.4]
  assign DualPortRAM_5_clock = clock; // @[transfer.scala 93:20:@199.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  value = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_516 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_518 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_520 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_522 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_524 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_526 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_528 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_530 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_532 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_534 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_536 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_538 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_540 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_542 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_544 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_546 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_548 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_550 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_552 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_554 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_556 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_558 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_560 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_562 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_564 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_566 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_568 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_570 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_572 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_574 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_576 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_578 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_580 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_582 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_584 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_586 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_588 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_590 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_592 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_594 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_596 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_598 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_600 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_602 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_604 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_606 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_608 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_610 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_612 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_614 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_616 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_618 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_620 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_622 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_624 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_626 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_628 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_630 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_632 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_634 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_636 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_638 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_640 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_642 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  value_1 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      value <= 8'h0;
    end else begin
      if (io_input_valid) begin
        if (_T_38) begin
          value <= 8'h0;
        end else begin
          value <= _T_41;
        end
      end
    end
    _T_516 <= io_input_valid;
    _T_518 <= _T_516;
    _T_520 <= _T_518;
    _T_522 <= _T_520;
    _T_524 <= _T_522;
    _T_526 <= _T_524;
    _T_528 <= _T_526;
    _T_530 <= _T_528;
    _T_532 <= _T_530;
    _T_534 <= _T_532;
    _T_536 <= _T_534;
    _T_538 <= _T_536;
    _T_540 <= _T_538;
    _T_542 <= _T_540;
    _T_544 <= _T_542;
    _T_546 <= _T_544;
    _T_548 <= _T_546;
    _T_550 <= _T_548;
    _T_552 <= _T_550;
    _T_554 <= _T_552;
    _T_556 <= _T_554;
    _T_558 <= _T_556;
    _T_560 <= _T_558;
    _T_562 <= _T_560;
    _T_564 <= _T_562;
    _T_566 <= _T_564;
    _T_568 <= _T_566;
    _T_570 <= _T_568;
    _T_572 <= _T_570;
    _T_574 <= _T_572;
    _T_576 <= _T_574;
    _T_578 <= _T_576;
    _T_580 <= _T_578;
    _T_582 <= _T_580;
    _T_584 <= _T_582;
    _T_586 <= _T_584;
    _T_588 <= _T_586;
    _T_590 <= _T_588;
    _T_592 <= _T_590;
    _T_594 <= _T_592;
    _T_596 <= _T_594;
    _T_598 <= _T_596;
    _T_600 <= _T_598;
    _T_602 <= _T_600;
    _T_604 <= _T_602;
    _T_606 <= _T_604;
    _T_608 <= _T_606;
    _T_610 <= _T_608;
    _T_612 <= _T_610;
    _T_614 <= _T_612;
    _T_616 <= _T_614;
    _T_618 <= _T_616;
    _T_620 <= _T_618;
    _T_622 <= _T_620;
    _T_624 <= _T_622;
    _T_626 <= _T_624;
    _T_628 <= _T_626;
    _T_630 <= _T_628;
    _T_632 <= _T_630;
    _T_634 <= _T_632;
    _T_636 <= _T_634;
    _T_638 <= _T_636;
    _T_640 <= _T_638;
    _T_642 <= _T_640;
    if (reset) begin
      value_1 <= 8'h0;
    end else begin
      if (io_out_valid) begin
        if (_T_646) begin
          value_1 <= 8'h0;
        end else begin
          value_1 <= _T_649;
        end
      end
    end
  end
endmodule
